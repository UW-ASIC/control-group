`default_nettype none

module aes_fsm ();

endmodule