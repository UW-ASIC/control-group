`default_nettype none

module req_queue ();

endmodule