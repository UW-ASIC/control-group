`default_nettype none

module ser_des ();

endmodule