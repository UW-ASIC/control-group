`default_nettype none

module sha_fsm ();

endmodule