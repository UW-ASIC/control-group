`default_nettype none

module scoreboard ();

endmodule